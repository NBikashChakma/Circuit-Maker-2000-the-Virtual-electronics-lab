CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 55 208 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89887e-315 0
0
13 Logic Switch~
5 61 158 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89887e-315 0
0
14 Logic Display~
6 573 358 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
43556 0
0
14 Logic Display~
6 682 155 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
43556 1
0
5 4011~
219 443 374 0 3 22
0 6 6 3
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
8157 0 0
2
43556 2
0
5 4011~
219 579 171 0 3 22
0 5 4 2
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
5572 0 0
2
43556 3
0
5 4011~
219 429 243 0 3 22
0 6 7 4
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
8901 0 0
2
43556 4
0
5 4011~
219 423 99 0 3 22
0 8 6 5
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
7361 0 0
2
43556 5
0
5 4011~
219 195 177 0 3 22
0 8 7 6
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
4747 0 0
2
43556 6
0
12
3 1 2 0 0 4224 0 6 4 0 0 3
606 171
682 171
682 173
3 1 3 0 0 4224 0 5 3 0 0 3
470 374
573 374
573 376
3 2 4 0 0 8320 0 7 6 0 0 4
456 243
497 243
497 180
555 180
3 1 5 0 0 8320 0 8 6 0 0 4
450 99
495 99
495 162
555 162
0 2 6 0 0 8192 0 0 5 6 0 3
343 365
343 383
419 383
0 1 6 0 0 4224 0 0 5 9 0 3
269 177
269 365
419 365
0 2 7 0 0 8320 0 0 7 11 0 3
131 186
131 252
405 252
0 1 8 0 0 8320 0 0 8 12 0 3
128 168
128 90
399 90
3 0 6 0 0 0 0 9 0 0 10 2
222 177
336 177
2 1 6 0 0 0 0 8 7 0 0 4
399 108
336 108
336 234
405 234
1 2 7 0 0 0 0 1 9 0 0 4
67 208
86 208
86 186
171 186
1 1 8 0 0 0 0 2 9 0 0 5
73 158
73 159
85 159
85 168
171 168
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
945 548 1062 572
955 556 1051 572
12 1  1   0   1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
953 494 1070 518
963 502 1059 518
12 1   0   1  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
961 440 1070 464
971 448 1059 464
11 0  1  1   0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
962 399 1063 423
972 407 1052 423
10 0  0  0  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
963 329 1080 353
973 337 1069 353
12 A  B    S  C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
646 346 707 370
656 354 696 370
5 carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
760 154 805 178
770 162 794 178
3 sum
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
