CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 117 131 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9196 0 0
2
43556.6 0
0
13 Logic Switch~
5 122 244 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3857 0 0
2
43556.6 1
0
13 Logic Switch~
5 124 184 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7125 0 0
2
43556.6 2
0
14 Logic Display~
6 660 292 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3641 0 0
2
43556.6 3
0
5 4071~
219 572 307 0 3 22
0 5 3 4
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
9821 0 0
2
43556.6 4
0
5 4081~
219 464 264 0 3 22
0 7 6 5
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
3187 0 0
2
43556.6 5
0
5 4081~
219 241 306 0 3 22
0 2 8 3
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
762 0 0
2
43556.6 6
0
14 Logic Display~
6 563 91 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
39 0 0
2
43556.6 7
0
5 4030~
219 442 105 0 3 22
0 7 6 9
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
9450 0 0
2
43556.6 8
0
5 4030~
219 234 166 0 3 22
0 2 8 7
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
3236 0 0
2
43556.6 9
0
12
1 1 2 0 0 4096 0 1 10 0 0 3
129 131
218 131
218 157
3 2 3 0 0 4224 0 7 5 0 0 3
262 306
559 306
559 316
1 3 4 0 0 8320 0 4 5 0 0 5
660 310
660 308
598 308
598 307
605 307
1 3 5 0 0 4224 0 5 6 0 0 4
559 298
516 298
516 264
485 264
0 2 6 0 0 8192 0 0 6 10 0 3
265 244
265 273
440 273
0 1 7 0 0 8320 0 0 6 11 0 3
311 165
311 255
440 255
0 2 8 0 0 4224 0 0 7 12 0 3
166 184
166 315
217 315
0 1 2 0 0 4224 0 0 7 1 0 3
188 131
188 297
217 297
3 1 9 0 0 8320 0 9 8 0 0 3
475 105
475 109
563 109
1 2 6 0 0 4224 0 2 9 0 0 4
134 244
409 244
409 114
426 114
1 3 7 0 0 0 0 9 10 0 0 6
426 96
368 96
368 165
270 165
270 166
267 166
1 2 8 0 0 0 0 3 10 0 0 4
136 184
214 184
214 175
218 175
13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
854 162 947 186
864 170 936 186
9 s   carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
849 216 1046 240
859 224 1035 240
22 A  B  Cin    S     Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
847 265 996 289
857 273 985 289
16 0  0  0    0   0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
855 322 996 346
865 330 985 346
15 0 0  1    1   0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
856 371 997 395
866 379 986 395
15 0  1  0   1   0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
861 436 1026 460
871 444 1015 460
18 0    1    1   0  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
837 502 954 526
847 510 943 526
12 1  0   0   1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
853 561 1002 585
863 569 991 585
16 1  0  1   0    1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
839 628 988 652
849 636 977 652
16 1  1   0   0   1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
834 723 967 747
844 731 956 747
14 1  1  1  1   1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1003 506 1032 530
1013 514 1021 530
1 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
593 84 622 108
603 92 611 108
1 s
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
669 323 714 347
679 331 703 347
3 Cin
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
