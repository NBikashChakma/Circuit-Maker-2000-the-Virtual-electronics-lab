CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 123 284 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
43556 0
0
13 Logic Switch~
5 118 249 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3472 0 0
2
43556 1
0
14 Logic Display~
6 698 138 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.89887e-315 0
0
14 Logic Display~
6 670 229 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
43556 2
0
9 2-In NOR~
219 558 246 0 3 22
0 4 6 5
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 0 0
1 U
4597 0 0
2
43556 3
0
9 2-In NOR~
219 373 158 0 3 22
0 8 7 4
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 0 0
1 U
3835 0 0
2
43556 4
0
9 2-In NOR~
219 226 358 0 3 22
0 2 2 7
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 0 0
1 U
3670 0 0
2
43556 5
0
9 2-In NOR~
219 217 258 0 3 22
0 3 2 6
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 0 0
1 U
5616 0 0
2
43556 6
0
9 2-In NOR~
219 215 163 0 3 22
0 3 3 8
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 0 0
1 U
9323 0 0
2
43556 7
0
16
0 0 2 0 0 4224 0 0 0 13 12 2
145 267
145 349
0 0 3 0 0 4224 0 0 0 14 16 2
140 249
140 154
1 0 4 0 0 4096 0 3 0 0 4 3
698 156
670 156
670 161
0 0 4 0 0 4224 0 0 0 7 0 3
412 161
670 161
670 157
1 0 3 0 0 0 0 2 0 0 14 2
130 249
130 249
3 1 5 0 0 4224 0 5 4 0 0 3
597 246
670 246
670 247
3 1 4 0 0 0 0 6 5 0 0 3
412 158
412 237
545 237
3 2 6 0 0 4224 0 8 5 0 0 4
256 258
534 258
534 255
545 255
3 2 7 0 0 8320 0 7 6 0 0 4
265 358
339 358
339 167
360 167
3 1 8 0 0 4224 0 9 6 0 0 4
254 163
339 163
339 149
360 149
0 2 2 0 0 0 0 0 7 12 0 3
176 349
176 367
213 367
0 1 2 0 0 0 0 0 7 0 0 3
138 350
138 349
213 349
1 2 2 0 0 0 0 1 8 0 0 4
135 284
134 284
134 267
204 267
0 1 3 0 0 0 0 0 8 0 0 3
127 250
127 249
204 249
0 2 3 0 0 0 0 0 9 16 0 3
162 154
162 172
202 172
0 1 3 0 0 0 0 0 9 0 0 3
128 153
128 154
202 154
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
923 235 1040 259
933 243 1029 259
12 A  B    S  C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
922 305 1023 329
932 313 1012 329
10 0  0  0  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
921 346 1030 370
931 354 1019 370
11 0  1  1   0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
913 400 1030 424
923 408 1019 424
12 1   0   1  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
905 454 1022 478
915 462 1011 478
12 1  1   0   1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
295 488 452 512
305 496 441 512
17 HALF ADDER TO NOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
74 274 103 298
84 282 92 298
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
62 235 91 259
72 243 80 259
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
761 133 822 157
771 141 811 157
5 carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
684 264 729 288
694 272 718 288
3 sum
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
