CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 48 225 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3835 0 0
2
43556.7 0
0
13 Logic Switch~
5 64 104 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3670 0 0
2
43556.7 0
0
14 Logic Display~
6 802 64 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5616 0 0
2
43556.7 0
0
5 4001~
219 700 82 0 3 22
0 4 4 3
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 2 0
1 U
9323 0 0
2
43556.7 0
0
5 4001~
219 485 56 0 3 22
0 5 6 4
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U1D
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 1 0
1 U
317 0 0
2
43556.7 0
0
5 4001~
219 363 172 0 3 22
0 5 7 6
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U1C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 1 0
1 U
3108 0 0
2
43556.7 0
0
5 4001~
219 190 234 0 3 22
0 8 8 7
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U1B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 1 0
1 U
4299 0 0
2
43556.7 0
0
5 4001~
219 183 102 0 3 22
0 2 2 5
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 1 0
1 U
9672 0 0
2
43556.7 0
0
13
1 0 2 0 0 0 0 2 0 0 13 2
76 104
76 104
3 1 3 0 0 4224 0 4 3 0 0 2
739 82
802 82
0 2 4 0 0 8192 0 0 4 4 0 3
654 73
654 91
687 91
3 1 4 0 0 12416 0 5 4 0 0 4
524 56
590 56
590 73
687 73
1 0 5 0 0 4224 0 5 0 0 9 3
472 47
308 47
308 163
3 2 6 0 0 8320 0 6 5 0 0 4
402 172
442 172
442 65
472 65
0 3 7 0 0 4096 0 0 7 8 0 3
261 181
261 234
229 234
2 0 7 0 0 4224 0 6 0 0 0 2
350 181
258 181
3 1 5 0 0 0 0 8 6 0 0 3
222 102
222 163
350 163
0 2 8 0 0 8192 0 0 7 11 0 3
112 225
112 243
177 243
1 1 8 0 0 4224 0 7 1 0 0 2
177 225
60 225
0 2 2 0 0 8320 0 0 8 13 0 3
112 104
112 111
170 111
1 0 2 0 0 128 0 8 0 0 0 4
170 93
112 93
112 104
73 104
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
