CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 156 430 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4459 0 0
2
43556.6 0
0
13 Logic Switch~
5 153 178 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3760 0 0
2
43556.6 1
0
14 Logic Display~
6 703 403 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
754 0 0
2
43556.6 2
0
14 Logic Display~
6 696 244 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9767 0 0
2
43556.6 3
0
5 4011~
219 625 420 0 3 22
0 6 6 4
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
7978 0 0
2
43556.6 4
0
5 4011~
219 611 263 0 3 22
0 7 6 5
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
3142 0 0
2
43556.6 5
0
5 4011~
219 431 422 0 3 22
0 8 2 6
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
3284 0 0
2
43556.6 6
0
5 4011~
219 408 187 0 3 22
0 3 8 7
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
659 0 0
2
43556.6 7
0
5 4011~
219 262 320 0 3 22
0 3 2 8
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
3800 0 0
2
43556.6 8
0
14
1 0 2 0 0 4096 0 1 0 0 11 2
168 430
168 431
1 0 3 0 0 4096 0 2 0 0 13 2
165 178
165 179
3 1 4 0 0 4224 0 5 3 0 0 3
652 420
703 420
703 421
3 1 5 0 0 4224 0 6 4 0 0 3
638 263
696 263
696 262
0 0 6 0 0 4096 0 0 0 8 6 2
493 422
557 422
1 2 6 0 0 0 0 5 5 0 0 4
601 411
557 411
557 429
601 429
3 1 7 0 0 8320 0 8 6 0 0 3
435 187
435 254
587 254
3 2 6 0 0 8320 0 7 6 0 0 4
458 422
493 422
493 272
587 272
3 0 8 0 0 4096 0 9 0 0 10 2
289 320
357 320
1 2 8 0 0 8320 0 7 8 0 0 4
407 413
357 413
357 196
384 196
0 0 2 0 0 4096 0 0 0 12 0 2
221 431
162 431
2 2 2 0 0 12416 0 9 7 0 0 4
238 329
221 329
221 431
407 431
0 0 3 0 0 4096 0 0 0 14 0 2
221 179
162 179
1 1 3 0 0 12416 0 9 8 0 0 4
238 311
221 311
221 178
384 178
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
731 239 760 263
741 247 749 263
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
766 428 803 452
776 436 792 452
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
918 137 1027 161
928 145 1016 161
11 TRUTH TABLE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
912 199 1037 223
922 207 1026 223
13 A  B   D   B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
926 260 1003 284
936 268 992 284
7 0 0 0 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
936 307 1013 331
946 315 1002 331
7 0 1 1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
931 363 1008 387
941 371 997 387
7 1 0 1 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
930 418 1007 442
940 426 996 442
7 1 1 0 0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
