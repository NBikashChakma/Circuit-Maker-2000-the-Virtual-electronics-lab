CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 31 125 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89887e-315 0
0
13 Logic Switch~
5 27 189 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
43640 0
0
13 Logic Switch~
5 43 339 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
43640 1
0
5 4001~
219 894 157 0 3 22
0 3 4 2
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 4 0
1 U
3421 0 0
2
43640 0
0
5 4001~
219 753 274 0 3 22
0 5 6 4
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U3D
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 3 0
1 U
8157 0 0
2
43640 0
0
5 4001~
219 630 151 0 3 22
0 7 6 5
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U3C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 3 0
1 U
5572 0 0
2
43640 0
0
5 4001~
219 428 51 0 3 22
0 10 8 7
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U3B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 3 0
1 U
8901 0 0
2
43640 0
0
5 4001~
219 766 31 0 3 22
0 7 5 3
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 3 0
1 U
7361 0 0
2
5.89887e-315 0
0
14 Logic Display~
6 972 37 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
43640 2
0
14 Logic Display~
6 1038 235 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
43640 3
0
5 4001~
219 905 317 0 3 22
0 4 6 11
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U2D
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 2 0
1 U
3472 0 0
2
43640 4
0
5 4001~
219 323 251 0 3 22
0 13 9 8
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U1C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 1 0
1 U
9998 0 0
2
43640 9
0
5 4001~
219 301 48 0 3 22
0 12 13 10
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U1B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 1 0
1 U
3536 0 0
2
43640 10
0
5 4001~
219 208 149 0 3 22
0 12 9 13
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 1 0
1 U
4597 0 0
2
43640 11
0
21
3 1 2 0 0 4224 0 4 9 0 0 4
933 157
933 65
972 65
972 55
1 3 3 0 0 8320 0 4 8 0 0 4
881 148
814 148
814 31
805 31
3 0 4 0 0 4096 0 5 0 0 4 2
792 274
857 274
1 2 4 0 0 8320 0 11 4 0 0 4
892 308
857 308
857 166
881 166
3 0 5 0 0 4096 0 6 0 0 15 2
669 151
730 151
0 2 6 0 0 4096 0 0 5 7 0 3
570 339
740 339
740 283
2 2 6 0 0 20608 0 6 11 0 0 8
617 160
570 160
570 339
391 339
391 399
879 399
879 326
892 326
1 0 7 0 0 8192 0 6 0 0 11 3
617 142
570 142
570 51
1 0 8 0 0 4224 0 3 0 0 12 3
55 339
391 339
391 251
0 0 9 0 0 4096 0 0 0 14 0 2
106 260
35 260
3 1 7 0 0 4224 0 7 8 0 0 6
467 51
684 51
684 0
743 0
743 22
753 22
2 3 8 0 0 0 0 7 12 0 0 4
415 60
391 60
391 251
362 251
3 1 10 0 0 4224 0 13 7 0 0 4
340 48
411 48
411 42
415 42
2 0 9 0 0 4224 0 12 0 0 20 3
310 260
106 260
106 156
1 2 5 0 0 8320 0 5 8 0 0 4
740 265
730 265
730 40
753 40
3 1 11 0 0 4224 0 11 10 0 0 3
944 317
1038 317
1038 253
0 1 12 0 0 8320 0 0 13 21 0 3
105 125
105 39
288 39
1 0 13 0 0 8192 0 12 0 0 19 3
310 242
252 242
252 150
2 3 13 0 0 8320 0 13 14 0 0 6
288 57
266 57
266 150
252 150
252 149
247 149
2 1 9 0 0 0 0 14 2 0 0 5
195 158
195 156
36 156
36 189
39 189
1 1 12 0 0 0 0 14 1 0 0 3
195 140
195 125
43 125
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
1612 325 1761 349
1622 333 1750 349
16 0  0  1   1    1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
1608 266 1749 290
1618 274 1738 290
15 0   0  0   0  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
1608 208 1757 232
1618 216 1746 232
16 A  B  Bi   D  B0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
