CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 101 222 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43556.5 0
0
13 Logic Switch~
5 85 167 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
43556.5 0
0
13 Logic Switch~
5 89 100 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
43556.5 0
0
5 4081~
219 764 334 0 3 22
0 4 3 5
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
3421 0 0
2
43556.5 0
0
5 4081~
219 426 268 0 3 22
0 10 6 2
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
8157 0 0
2
43556.5 0
0
14 Logic Display~
6 744 142 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
43556.5 0
0
14 Logic Display~
6 988 216 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
43556.5 0
0
5 4071~
219 879 267 0 3 22
0 2 5 8
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
7361 0 0
2
43556.5 0
0
5 4049~
219 576 297 0 2 22
0 9 4
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 2 0
1 U
4747 0 0
2
43556.5 0
0
5 4049~
219 263 256 0 2 22
0 11 10
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 2 0
1 U
972 0 0
2
43556.5 0
0
5 4030~
219 583 158 0 3 22
0 9 3 7
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
3472 0 0
2
43556.5 0
0
5 4030~
219 261 158 0 3 22
0 11 6 9
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
9998 0 0
2
43556.5 0
0
22
3 0 2 0 0 0 0 5 0 0 10 2
447 268
447 268
2 0 3 0 0 8192 0 4 0 0 13 3
740 343
740 342
711 342
1 0 4 0 0 8192 0 4 0 0 12 3
740 325
740 324
711 324
3 2 5 0 0 8320 0 4 8 0 0 3
785 334
785 276
866 276
1 0 3 0 0 0 0 1 0 0 15 2
113 222
113 221
1 0 6 0 0 0 0 2 0 0 8 2
97 167
97 167
1 0 7 0 0 4096 0 6 0 0 11 2
744 160
744 158
0 0 6 0 0 4096 0 0 0 21 0 2
139 167
86 167
3 1 8 0 0 4224 0 8 7 0 0 3
912 267
988 267
988 234
0 1 2 0 0 4224 0 0 8 0 0 4
443 268
816 268
816 258
866 258
3 0 7 0 0 4224 0 11 0 0 0 2
616 158
748 158
2 0 4 0 0 4224 0 9 0 0 0 4
597 297
681 297
681 324
720 324
0 0 3 0 0 8192 0 0 0 15 0 3
472 167
472 342
720 342
0 1 9 0 0 4096 0 0 9 16 0 3
516 149
516 297
561 297
2 0 3 0 0 4224 0 11 0 0 0 6
567 167
312 167
312 189
131 189
131 221
109 221
3 1 9 0 0 4224 0 12 11 0 0 4
294 158
455 158
455 149
567 149
2 0 6 0 0 4224 0 5 0 0 21 3
402 277
157 277
157 167
1 2 10 0 0 12416 0 5 10 0 0 4
402 259
392 259
392 256
284 256
0 0 11 0 0 4224 0 0 0 20 22 2
203 256
203 135
1 0 11 0 0 0 0 10 0 0 0 2
248 256
197 256
2 0 6 0 0 0 0 12 0 0 0 2
245 167
136 167
1 1 11 0 0 128 0 3 12 0 0 6
101 100
101 99
139 99
139 135
245 135
245 149
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
