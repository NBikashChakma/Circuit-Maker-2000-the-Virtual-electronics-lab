CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
250 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 89 409 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3649 0 0
2
43556.6 0
0
13 Logic Switch~
5 120 336 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3716 0 0
2
43556.6 1
0
13 Logic Switch~
5 126 164 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4797 0 0
2
43556.6 2
0
9 2-In NOR~
219 911 480 0 3 22
0 4 3 2
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4681 0 0
2
43556.6 3
0
14 Logic Display~
6 990 463 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9730 0 0
2
43556.6 4
0
14 Logic Display~
6 1118 231 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9874 0 0
2
43556.6 5
0
9 2-In NOR~
219 877 154 0 3 22
0 10 3 9
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 0 0
1 U
364 0 0
2
43556.6 6
0
9 2-In NOR~
219 1008 247 0 3 22
0 9 8 7
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U2D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3656 0 0
2
43556.6 7
0
9 2-In NOR~
219 874 346 0 3 22
0 3 5 8
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U2C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3131 0 0
2
43556.6 8
0
9 2-In NOR~
219 679 254 0 3 22
0 10 5 3
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6772 0 0
2
43556.6 9
0
9 2-In NOR~
219 531 248 0 3 22
0 11 12 10
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
9557 0 0
2
43556.6 10
0
9 2-In NOR~
219 370 328 0 3 22
0 4 13 12
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
5789 0 0
2
43556.6 11
0
9 2-In NOR~
219 379 172 0 3 22
0 6 4 11
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7328 0 0
2
43556.6 12
0
9 2-In NOR~
219 210 241 0 3 22
0 6 13 4
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4799 0 0
2
43556.6 13
0
22
3 1 2 0 0 4224 0 4 5 0 0 3
950 480
990 480
990 481
0 2 3 0 0 4224 0 0 4 10 0 5
775 254
775 496
872 496
872 489
898 489
0 1 4 0 0 8320 0 0 4 21 0 5
282 241
282 460
865 460
865 471
898 471
1 0 5 0 0 4096 0 1 0 0 14 2
101 409
101 408
1 0 6 0 0 4096 0 3 0 0 20 2
138 164
138 163
3 1 7 0 0 4224 0 8 6 0 0 3
1047 247
1118 247
1118 249
3 2 8 0 0 4224 0 9 8 0 0 3
913 346
913 256
995 256
3 1 9 0 0 4224 0 7 8 0 0 3
916 154
916 238
995 238
0 2 3 0 0 0 0 0 7 10 0 3
831 254
831 163
864 163
3 1 3 0 0 0 0 10 9 0 0 6
718 254
831 254
831 340
846 340
846 337
861 337
0 2 5 0 0 12288 0 0 9 14 0 4
636 308
719 308
719 355
861 355
0 1 10 0 0 8320 0 0 7 13 0 3
629 248
629 145
864 145
1 3 10 0 0 0 0 10 11 0 0 3
666 245
666 248
570 248
2 0 5 0 0 12416 0 10 0 0 0 4
666 263
636 263
636 408
97 408
3 1 11 0 0 4224 0 13 11 0 0 4
418 172
491 172
491 239
518 239
3 2 12 0 0 4224 0 12 11 0 0 4
409 328
491 328
491 257
518 257
2 0 13 0 0 8192 0 14 0 0 19 3
197 250
164 250
164 337
1 0 6 0 0 8192 0 14 0 0 20 3
197 232
164 232
164 163
2 1 13 0 0 4224 0 12 2 0 0 3
357 337
132 337
132 336
1 0 6 0 0 4224 0 13 0 0 0 2
366 163
134 163
3 0 4 0 0 0 0 14 0 0 22 2
249 241
315 241
1 2 4 0 0 0 0 12 13 0 0 4
357 319
315 319
315 181
366 181
13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
957 500 986 524
967 508 975 524
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
135 422 196 446
145 430 185 446
5 carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1146 239 1191 263
1156 247 1180 263
3 sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
1442 196 1583 220
1452 204 1572 220
15 A  B  C   S   C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
1434 239 1583 263
1444 247 1572 263
16 0    0   0  0  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1428 276 1553 300
1438 284 1542 300
13 0    0   1  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1553 280 1582 304
1563 288 1571 304
1 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1443 322 1568 346
1453 330 1557 346
13 0 1  1   0  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1432 374 1557 398
1442 382 1546 398
13 1  0  0  1  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
1424 421 1557 445
1434 429 1546 445
14 1  0  1   0  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
1431 465 1564 489
1441 473 1553 489
14 1  1  0   0  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
1420 509 1553 533
1430 517 1542 533
14 1  1 1   1   1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1590 308 1707 332
1600 316 1696 332
12 0 1 0   1  0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
