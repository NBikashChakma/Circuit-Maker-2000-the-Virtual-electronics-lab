CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 24 493 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7168 0 0
2
43556.6 0
0
13 Logic Switch~
5 28 425 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
631 0 0
2
43556.6 1
0
13 Logic Switch~
5 27 115 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9466 0 0
2
43556.6 2
0
14 Logic Display~
6 976 494 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3266 0 0
2
43556.6 3
0
14 Logic Display~
6 940 285 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7693 0 0
2
43556.6 4
0
5 4011~
219 888 526 0 3 22
0 8 7 5
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
3723 0 0
2
43556.6 5
0
5 4011~
219 875 303 0 3 22
0 9 8 6
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
3440 0 0
2
43556.6 6
0
5 4011~
219 733 483 0 3 22
0 11 2 8
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
6263 0 0
2
43556.6 7
0
5 4011~
219 708 248 0 3 22
0 10 11 9
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
4900 0 0
2
43556.6 8
0
5 4011~
219 575 340 0 3 22
0 10 2 11
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
8783 0 0
2
43556.6 9
0
5 4011~
219 461 238 0 3 22
0 12 7 10
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
3221 0 0
2
43556.6 10
0
5 4011~
219 334 417 0 3 22
0 13 3 7
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
3215 0 0
2
43556.6 11
0
5 4011~
219 311 125 0 3 22
0 4 13 12
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
7903 0 0
2
43556.6 12
0
5 4011~
219 158 290 0 3 22
0 4 3 13
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
7121 0 0
2
43556.6 13
0
23
1 0 2 0 0 4096 0 1 0 0 12 2
36 493
36 492
1 0 3 0 0 4096 0 2 0 0 22 2
40 425
40 426
1 0 4 0 0 4096 0 3 0 0 23 2
39 115
39 116
3 1 5 0 0 8320 0 6 4 0 0 4
915 526
915 541
976 541
976 512
3 1 6 0 0 4224 0 7 5 0 0 2
902 303
940 303
2 3 7 0 0 4224 0 6 12 0 0 7
864 535
358 535
358 502
375 502
375 483
361 483
361 417
0 1 8 0 0 8192 0 0 6 8 0 3
784 483
784 517
864 517
3 2 8 0 0 8320 0 8 7 0 0 4
760 483
800 483
800 312
851 312
3 1 9 0 0 12416 0 9 7 0 0 4
735 248
766 248
766 294
851 294
2 0 2 0 0 8192 0 10 0 0 12 3
551 349
529 349
529 492
1 0 10 0 0 8192 0 10 0 0 15 3
551 331
529 331
529 238
2 0 2 0 0 4224 0 8 0 0 0 2
709 492
31 492
3 0 11 0 0 4096 0 10 0 0 14 2
602 340
644 340
2 1 11 0 0 8320 0 9 8 0 0 4
684 257
644 257
644 474
709 474
3 1 10 0 0 4224 0 11 9 0 0 3
488 238
684 238
684 239
2 3 7 0 0 0 0 11 12 0 0 6
437 247
360 247
360 380
376 380
376 417
361 417
3 1 12 0 0 8320 0 13 11 0 0 4
338 125
362 125
362 229
437 229
3 0 13 0 0 4096 0 14 0 0 19 2
185 290
255 290
2 1 13 0 0 8320 0 13 12 0 0 4
287 134
255 134
255 408
310 408
1 0 4 0 0 8192 0 14 0 0 23 3
134 281
110 281
110 116
2 0 3 0 0 8192 0 14 0 0 22 3
134 299
110 299
110 426
2 0 3 0 0 4224 0 12 0 0 0 2
310 426
34 426
1 0 4 0 0 4224 0 13 0 0 0 2
287 116
32 116
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1011 550 1048 574
1021 558 1037 574
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
982 285 1011 309
992 293 1000 309
1 D
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
