CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 137 504 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6901 0 0
2
43556.7 0
0
13 Logic Switch~
5 81 327 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
842 0 0
2
5.89887e-315 0
0
13 Logic Switch~
5 87 281 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3277 0 0
2
5.89887e-315 5.26354e-315
0
14 Logic Display~
6 1171 553 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
43556.7 1
0
14 Logic Display~
6 1340 340 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
5.89887e-315 5.30499e-315
0
5 4011~
219 1229 359 0 3 22
0 7 8 6
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
5551 0 0
2
5.89887e-315 5.32571e-315
0
5 4011~
219 834 570 0 3 22
0 10 2 9
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
6986 0 0
2
5.89887e-315 5.34643e-315
0
5 4011~
219 892 495 0 3 22
0 10 3 8
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
8745 0 0
2
5.89887e-315 5.3568e-315
0
5 4011~
219 878 277 0 3 22
0 11 10 7
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
9592 0 0
2
5.89887e-315 5.36716e-315
0
5 4011~
219 732 391 0 3 22
0 11 3 10
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
8748 0 0
2
5.89887e-315 5.37752e-315
0
5 4011~
219 569 268 0 3 22
0 13 12 11
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
7168 0 0
2
5.89887e-315 5.38788e-315
0
5 4011~
219 368 420 0 3 22
0 2 4 12
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
631 0 0
2
5.89887e-315 5.39306e-315
0
5 4011~
219 351 122 0 3 22
0 5 2 13
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
9466 0 0
2
5.89887e-315 5.39824e-315
0
5 4011~
219 185 290 0 3 22
0 5 4 2
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 0 0
1 U
3266 0 0
2
5.89887e-315 5.40342e-315
0
23
2 0 2 0 0 4224 0 7 0 0 18 3
810 579
226 579
226 290
1 0 3 0 0 0 0 1 0 0 11 2
149 504
149 504
1 0 4 0 0 4096 0 2 0 0 22 2
93 327
93 326
1 0 5 0 0 0 0 3 0 0 23 2
99 281
99 281
3 1 6 0 0 4224 0 6 5 0 0 3
1256 359
1340 359
1340 358
3 1 7 0 0 4224 0 9 6 0 0 4
905 277
1144 277
1144 350
1205 350
3 2 8 0 0 4224 0 8 6 0 0 4
919 495
1149 495
1149 368
1205 368
3 1 9 0 0 4224 0 7 4 0 0 3
861 570
1171 570
1171 571
0 1 10 0 0 4096 0 0 7 12 0 3
781 391
781 561
810 561
2 0 3 0 0 8192 0 10 0 0 11 3
708 400
662 400
662 504
2 0 3 0 0 4224 0 8 0 0 0 2
868 504
144 504
3 0 10 0 0 0 0 10 0 0 13 2
759 391
845 391
1 2 10 0 0 8320 0 8 9 0 0 4
868 486
845 486
845 286
854 286
0 1 11 0 0 4224 0 0 9 15 0 2
661 268
854 268
3 1 11 0 0 0 0 11 10 0 0 4
596 268
661 268
661 382
708 382
3 2 12 0 0 8320 0 12 11 0 0 3
395 420
395 277
545 277
3 1 13 0 0 8320 0 13 11 0 0 3
378 122
378 259
545 259
3 0 2 0 0 0 0 14 0 0 21 2
212 290
265 290
0 1 5 0 0 8320 0 0 13 23 0 3
143 281
143 113
327 113
2 0 4 0 0 4224 0 12 0 0 22 3
344 429
143 429
143 299
2 1 2 0 0 0 0 13 12 0 0 4
327 131
265 131
265 411
344 411
0 2 4 0 0 0 0 0 14 0 0 4
89 326
102 326
102 299
161 299
0 1 5 0 0 0 0 0 14 0 0 2
96 281
161 281
18
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1232 87 1280 110
1245 97 1266 112
3 1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1239 124 1285 147
1251 134 1272 149
3 2 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
1107 684 1253 707
1120 694 1239 709
17 C = A.B+Ci(A(+)B)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
975 122 1084 145
987 132 1071 147
12 S=A(+)B(+)Ci
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
175 1405 270 1428
187 1415 257 1430
10 1 1 1 1  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
162 1357 273 1380
175 1367 259 1382
12 1 1  0  0  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
170 1302 279 1325
182 1312 266 1327
12 1 0  1  0  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
170 1232 286 1255
182 1242 273 1257
13 1  0  0   1 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
182 1167 300 1190
195 1177 286 1192
13 0  1  1  0  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
186 1114 297 1137
199 1124 283 1139
12 0  1 0  1  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
196 1041 314 1064
209 1051 300 1066
13 0  0  1  1  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
200 956 330 979
212 966 317 981
15 0  0  0   0   0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
199 885 372 908
211 895 359 910
21 A   B   Ci     S    C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
104 501 141 525
114 509 130 525
2 ci
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
43 262 72 286
53 270 61 286
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
42 339 71 363
52 347 60 363
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1385 311 1418 334
1397 321 1405 336
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1221 567 1256 590
1234 577 1242 592
1 C
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
