CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 150 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
7
13 Logic Switch~
5 127 283 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4212 0 0
2
43556.6 0
0
13 Logic Switch~
5 125 205 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4720 0 0
2
43556.6 1
0
13 Logic Switch~
5 115 107 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5551 0 0
2
43556.6 2
0
14 Logic Display~
6 605 155 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6986 0 0
2
43556.6 3
0
5 4071~
219 541 171 0 3 22
0 7 6 5
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
8745 0 0
2
43556.6 4
0
5 4081~
219 405 247 0 3 22
0 3 2 6
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
9592 0 0
2
43556.6 5
0
5 4049~
219 227 139 0 2 22
0 4 7
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U1A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
8748 0 0
2
43556.6 6
0
13
1 0 2 0 0 0 0 1 0 0 10 2
139 283
139 283
1 0 3 0 0 0 0 2 0 0 11 2
137 205
137 205
1 0 4 0 0 0 0 3 0 0 13 2
127 107
127 107
1 0 5 0 0 4096 0 4 0 0 5 2
605 173
605 171
3 0 5 0 0 4224 0 5 0 0 0 2
574 171
611 171
2 0 6 0 0 4096 0 5 0 0 0 2
528 180
535 180
3 2 6 0 0 8320 0 6 5 0 0 4
426 247
483 247
483 180
528 180
2 1 7 0 0 4224 0 7 5 0 0 4
248 139
483 139
483 162
528 162
1 0 4 0 0 4096 0 7 0 0 12 2
212 139
212 140
0 2 2 0 0 4224 0 0 6 0 0 4
134 283
295 283
295 256
381 256
0 1 3 0 0 4224 0 0 6 0 0 4
133 205
295 205
295 238
381 238
0 0 4 0 0 4096 0 0 0 13 0 3
189 107
189 140
217 140
0 0 4 0 0 4224 0 0 0 0 0 2
123 107
296 107
16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
842 748 967 772
852 756 956 772
13 1   1   1   1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
848 698 957 722
858 706 946 722
11 1  1  0   0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
844 635 953 659
854 643 942 659
11 1  0  1   0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
863 556 964 580
873 564 953 580
10 1  0  0  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
861 503 970 527
871 511 959 527
11 0   1  1  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
854 449 955 473
864 457 944 473
10 0  1  0  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
869 394 970 418
879 402 959 418
10 0  0  1  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
866 323 967 347
876 331 956 347
10 0  0  0  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
875 266 1000 290
885 274 989 290
13 p  q   r    y
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
594 191 679 215
604 199 668 215
8 S=P*+Q.R
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
568 135 597 159
578 143 586 159
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
436 249 481 273
446 257 470 273
3 Q.R
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
153 257 182 281
163 265 171 281
1 R
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
145 174 174 198
155 182 163 198
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
123 76 152 100
133 84 141 100
1 p
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
245 143 282 167
255 151 271 167
2 P*
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
